module dataPath(/*INPUTS GO HERE*/);

endmodule // dataPath
